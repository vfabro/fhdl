architecture a of myEntity is
begin
  process 
  begin
   a <= myFunction (c);
  end process;
end architecture;
