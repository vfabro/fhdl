architecture x of myEntity is
begin 
  a <= mySignal (a'high downto a'low);
  c <= mySignal (x'attrDesignator);
end;
